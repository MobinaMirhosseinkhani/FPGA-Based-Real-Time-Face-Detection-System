module dense_layer(
    input clk,
    input rst, 
    output reg out
);
    reg [31:0] weights [0:199];  // ????? ????? ????? ???? ??????
    reg [31:0] bias [0:1];
    integer i, j;
    reg [1:0] output_data;
    reg [1:0] temp_output; 
    reg [31:0] input_data [99:0];

initial
begin
	bias[0]=32'h3F27D4FE;
	bias[01]=32'h3F27D4FE;
		
weights[0]=32'hBEC1C283;
weights[1]=32'h3F0A4075;
weights[2]=32'h3F2DCB21;
weights[3]=32'hBE7AEAE0;
weights[4]=32'hBE692930;
weights[5]=32'h3D8551E4;
weights[6]=32'hBF40A5F6;
weights[7]=32'h3F2CDBF5;
weights[8]=32'hBF173B19;
weights[9]=32'h3F5793D7;
weights[10]=32'hBF4B2135;
weights[11]=32'h3F1EAAA3;
weights[12]=32'hBF402620;
weights[13]=32'h3F822F5C;
weights[14]=32'hBF16B54D;
weights[15]=32'h3F471755;
weights[16]=32'h3EA69AC8;
weights[17]=32'hBEAF9F0F;
weights[18]=32'hBE8FA82D;
weights[19]=32'h3E0BC16B;
weights[20]=32'hBF33260F;
weights[21]=32'h3F04F23B;
weights[22]=32'hBEB9442A;
weights[23]=32'h3DF124AD;
weights[24]=32'hBFB24F3E;
weights[25]=32'h3FB74434;
weights[26]=32'h3E9F553C;
weights[27]=32'hBE02D423;
weights[28]=32'hBDE495F1;
weights[29]=32'h3DCD3BAB;
weights[30]=32'hBDF8211C;
weights[31]=32'hBE90889B;
weights[32]=32'hBEA46777;
weights[33]=32'h3EB46872;
weights[34]=32'hBFA6109E;
weights[35]=32'h3FAB1CD2;
weights[36]=32'hBF340694;
weights[37]=32'h3F523178;
weights[38]=32'hBD7F5599;
weights[39]=32'h3E57B7F8;
weights[40]=32'h3E4E2D81;
weights[41]=32'h3E314E46;
weights[42]=32'hBFEEECA0;
weights[43]=32'h4007FD5E;
weights[44]=32'hBF2FE4B0;
weights[45]=32'h3EF40AF6;
weights[46]=32'h3F1FAC8D;
weights[47]=32'hBF42E7DC;
weights[48]=32'h3F230C1C;
weights[49]=32'hBF44B6F8;
weights[50]=32'h3F5610ED;
weights[51]=32'hBF1A97AB;
weights[52]=32'h3F3AFD1F;
weights[53]=32'hBF459DC5;
weights[54]=32'hBF0833CA;
weights[55]=32'h3F2D6978;
weights[56]=32'hBFEF5245;
weights[57]=32'h3FF5EABD;
weights[58]=32'h3E7E26B7;
weights[59]=32'hBDDD44E3;
weights[60]=32'hBD90AECF;
weights[61]=32'h3EC6C066;
weights[62]=32'h3FD16960;
weights[63]=32'hBF9618DA;
weights[64]=32'hBD5D3183;
weights[65]=32'h3DDF943A;
weights[66]=32'h3F176A60;
weights[67]=32'hBF2F7802;
weights[68]=32'h3FFB236A;
weights[69]=32'hC00E7D24;
weights[70]=32'h401DBAD4;
weights[71]=32'hC01C3D8E;
weights[72]=32'h3EDF8C33;
weights[73]=32'hBF1CD14B;
weights[74]=32'h3DDE385B;
weights[75]=32'hBE077AB4;
weights[76]=32'h3F8C51A8;
weights[77]=32'hBF7857BA;
weights[78]=32'hBF01B24E;
weights[79]=32'h3F15DA66;
weights[80]=32'h3E3875CA;
weights[81]=32'h3DBC088F;
weights[82]=32'hBED49BC6;
weights[83]=32'hBD37F41E;
weights[84]=32'hBD50B006;
weights[85]=32'h3D99DB51;
weights[86]=32'h3EFD2E40;
weights[87]=32'hBEF628D9;
weights[88]=32'h3F5483DC; 
weights[89]=32'hBF492646;
weights[90]=32'h3FA98500;
weights[91]=32'hBFBD2B7F;
weights[92]=32'h3F9150AA;
weights[93]=32'hBF87E17B;
weights[94]=32'h3DAAB1DD;
weights[95]=32'hBDA7AD16;
weights[96]=32'hBE064DD4;
weights[97]=32'h3E85AE55;
weights[98]=32'hBF00D8B6;
weights[99]=32'h3F0D318E;
weights[100]=32'hBECA7DF3;
weights[101]=32'h3EC33B84;
weights[102]=32'hBE7B8C0F;
weights[103]=32'h3E88C10A;
weights[104]=32'h3F7B38D9;
weights[105]=32'hBF828C3E;
weights[106]=32'h3FBE065C;
weights[107]=32'hBFDCE51D;
weights[108]=32'hBF9C525C;
weights[109]=32'h3F56A17B;
weights[110]=32'hBF1C109C;
weights[111]=32'h3F201278;
weights[112]=32'h3FEC9FC1;
weights[113]=32'hBFE23B4E;
weights[114]=32'h3F9B3401;
weights[115]=32'hBF757CB3;
weights[116]=32'hBEFB8839;
weights[117]=32'h3E83D018;
weights[118]=32'hBF3F7041;
weights[119]=32'h3F27B431;
weights[120]=32'hBE0204AE;
weights[121]=32'h3D570233;
weights[122]=32'hBD205199;
weights[123]=32'h3D000ECA;
weights[124]=32'hBD4B36E1;
weights[125]=32'h3D2746B9;
weights[126]=32'hBB4091A8;
weights[127]=32'hBE929034;
weights[128]=32'hBEAB4C61;
weights[129]=32'h3EE59AA3;
weights[130]=32'h3D6B985A;
weights[131]=32'h3B8635E1;
weights[132]=32'hBE876B6C;
weights[133]=32'h3E10E57F;
weights[134]=32'h3EB3D059;
weights[135]=32'hBE4FAD84;
weights[136]=32'hBE544F4E;
weights[137]=32'h3F0835DC;
weights[138]=32'hBF00F6F9;
weights[139]=32'h3EF550FB;
weights[140]=32'h3EDDBCF3;
weights[141]=32'hBE77027B;
weights[142]=32'hBF1DC0B6;
weights[143]=32'h3F5A4A51;
weights[144]=32'hBE2A9AC8;
weights[145]=32'hBE08EC36;
weights[146]=32'h3E73EF03;
weights[147]=32'hBE15D165;
weights[148]=32'h3EDDDD38;
weights[149]=32'hBF2F6215;
weights[150]=32'h3F255959;
weights[151]=32'hBF20F2F9;
weights[152]=32'h3E786FC4;
weights[153]=32'hBE060FC3;
weights[154]=32'h3D646F0A;
weights[155]=32'hBEB1F8BE;
weights[156]=32'hBFBA3AC9;
weights[157]=32'h3FB4F38D;
weights[158]=32'h3EFDAAF5;
weights[159]=32'hBF39E21B;
weights[160]=32'h3F0E9B22;
weights[161]=32'hBF450DF4;
weights[162]=32'hBEDB025C;
weights[163]=32'h3EDADDE5;
weights[164]=32'hBEB33807;
weights[165]=32'h3EA34BE4;
weights[166]=32'hBF5B9067;
weights[167]=32'h3F631C5D;
weights[168]=32'h3EDB5F56;
weights[169]=32'hBE799BCE;
weights[170]=32'h3E1602C3;
weights[171]=32'hBEAD9164;
weights[172]=32'hBE864F6B;
weights[173]=32'h3F12E2A8;
weights[174]=32'hBED63690;
weights[175]=32'h3E7B8431;
weights[176]=32'hBF2307DE;
weights[177]=32'h3EB2AC08;
weights[178]=32'h3F7DB796;
weights[179]=32'hBF6CBA60;
weights[180]=32'h3F52CD77;
weights[181]=32'hBEF140A8;
weights[182]=32'hBD105A99;
weights[183]=32'hBEBC3061;
weights[184]=32'h3D9CCE46;
weights[185]=32'hBEA29097;
weights[186]=32'hBDAF4F91;
weights[187]=32'h3E231B55;
weights[188]=32'h3E657DCA;
weights[189]=32'h3DB23AF9;
weights[190]=32'h3D494B4B;
weights[191]=32'h3DFC2B9D;
weights[192]=32'h3DABEE9A;
weights[193]=32'hBDDB0068;
weights[194]=32'hBED60052;
weights[195]=32'h3D840676;
weights[196]=32'hBE904A05;
weights[197]=32'h3F05D4F2;
weights[198]=32'h3E7D961F;
weights[199]=32'hBEE769BE;


input_data[0] = 32'h9E ; 
input_data[1] = 32'h54 ; 
input_data[2] = 32'h8D ; 
input_data[3] = 32'h58 ; 
input_data[4] = 32'h58 ; 
input_data[5] = 32'h53 ; 
input_data[6] = 32'h59 ; 
input_data[7] = 32'h5A ; 
input_data[8] = 32'h2D ; 
input_data[9] = 32'hA9 ; 
input_data[10] = 32'hA7 ; 
input_data[11] = 32'h58 ; 
input_data[12] = 32'hA9 ; 
input_data[13] = 32'h63 ; 
input_data[14] = 32'h5C ; 
input_data[15] = 32'h54 ; 
input_data[16] = 32'h5D ; 
input_data[17] = 32'h5C ; 
input_data[18] = 32'h34 ; 
input_data[19] = 32'hB4 ; 
input_data[20] = 32'hAB ; 
input_data[21] = 32'hA2 ; 
input_data[22] = 32'h8A ; 
input_data[23] = 32'h26 ; 
input_data[24] = 32'h4B ; 
input_data[25] = 32'h59 ; 
input_data[26] = 32'h2E ; 
input_data[27] = 32'h2E ; 
input_data[28] = 32'h43 ; 
input_data[29] = 32'hBF ; 
input_data[30] = 32'hAE ; 
input_data[31] = 32'h7D ; 
input_data[32] = 32'h7D ; 
input_data[33] = 32'h37 ; 
input_data[34] = 32'h42 ; 
input_data[35] = 32'h37 ; 
input_data[36] = 32'h4F ; 
input_data[37] = 32'h32 ; 
input_data[38] = 32'h3B ; 
input_data[39] = 32'hC0 ; 
input_data[40] = 32'hAC ; 
input_data[41] = 32'hAE ; 
input_data[42] = 32'h8F ; 
input_data[43] = 32'h4A ; 
input_data[44] = 32'hB1 ; 
input_data[45] = 32'h55 ; 
input_data[46] = 32'h4C ; 
input_data[47] = 32'h5F ; 
input_data[48] = 32'h63 ; 
input_data[49] = 32'hC5 ; 
input_data[50] = 32'hAF ; 
input_data[51] = 32'hAD ; 
input_data[52] = 32'h9B ; 
input_data[53] = 32'h59 ; 
input_data[54] = 32'hC3 ; 
input_data[55] = 32'h68 ; 
input_data[56] = 32'h5F ; 
input_data[57] = 32'h5F ; 
input_data[58] = 32'hB3 ; 
input_data[59] = 32'hC5 ; 
input_data[60] = 32'hA6 ; 
input_data[61] = 32'h88 ; 
input_data[62] = 32'h67 ; 
input_data[63] = 32'h84 ; 
input_data[64] = 32'h58 ; 
input_data[65] = 32'h3B ; 
input_data[66] = 32'h53 ; 
input_data[67] = 32'h4B ; 
input_data[68] = 32'h7D ; 
input_data[69] = 32'h87 ; 
input_data[70] = 32'h76 ; 
input_data[71] = 32'h44 ; 
input_data[72] = 32'h41 ; 
input_data[73] = 32'h46 ; 
input_data[74] = 32'h3C ; 
input_data[75] = 32'h3E ; 
input_data[76] = 32'h42 ; 
input_data[77] = 32'h25 ; 
input_data[78] = 32'h7A ; 
input_data[79] = 32'h6F ; 
input_data[80] = 32'h6A ; 
input_data[81] = 32'h3B ; 
input_data[82] = 32'h33 ; 
input_data[83] = 32'h59 ; 
input_data[84] = 32'h32 ; 
input_data[85] = 32'h34 ; 
input_data[86] = 32'h2B ; 
input_data[87] = 32'h1D ; 
input_data[88] = 32'h74 ; 
input_data[89] = 32'h6F ; 
input_data[90] = 32'h63 ; 
input_data[91] = 32'h64 ; 
input_data[92] = 32'h20 ; 
input_data[93] = 32'h33 ; 
input_data[94] = 32'h1D ; 
input_data[95] = 32'h1E ; 
input_data[96] = 32'h39 ; 
input_data[97] = 32'h1F ; 
input_data[98] = 32'h6D ; 
input_data[99] = 32'h6C ;



end
 
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            output_data[0] <= 0;
            output_data[1] <= 0;
        end else begin
            for (j = 0; j < 2; j = j + 1) begin
                temp_output[j] = bias[j]; 
                for (i = 0; i < 100; i = i + 1) begin
                    temp_output[j] = temp_output[j] + (input_data[i] * weights[i+j*100]);
                end
            end
            
        
            output_data[0] <= temp_output[0];
            output_data[1] <= temp_output[1];
				 
			        if (output_data[0] > output_data[1])
            out <= 1'b0;
        else
            out <= 1'b1;
        end
        

    end
endmodule
